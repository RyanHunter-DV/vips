`ifndef Axi4MasterAgent__svh
`define Axi4MasterAgent__svh
`endif