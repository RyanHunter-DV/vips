`ifndef ChiVipIf__sv
`define ChiVipIf__sv

interface ChiVipIf#(REQCHN=1,RSPCHN=1,DATCHN=1,SNPCHN=1)(input clk,input resetn);
	


endinterface

`endif