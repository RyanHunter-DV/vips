`ifndef RhQLpiEnv__sv
`define RhQLpiEnv__sv

package RhQLpiEnv;

	import uvm_pkg::*;
	import RhLpiVip::*;

	`include "RhQLpiScoreboard.svh" 
	`include "RhQLpiEnv.svh"

endpackage

`endif