`ifndef Axi4SeqrBase__svh
`define Axi4SeqrBase__svh
`endif