`ifndef rh_axi4_ifcontrol_base__svh
`define rh_axi4_ifcontrol_base__svh

virtual class rh_axi4_ifcontrol_base;

    pure virtual function rh_axi4_vip_configBase createConfig(string name="cfg");

endclass


`endif
