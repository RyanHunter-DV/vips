`ifndef Axi4AgentBase__svh
`define Axi4AgentBase__svh
`endif