`ifndef Axi4Types__svh
`define Axi4Types__svh
`endif