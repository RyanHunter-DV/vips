`ifndef rh_ahbResetTrans__svh
`define rh_ahbResetTrans__svh

class rh_ahbResetTrans extends uvm_sequence_item; // {

	rh_resetAction_enum action;


endclass // }


`endif
