`ifndef rhaxi4_testBase__svh
`define rhaxi4_testBase__svh

class rhaxi4_testBase extends uvm_test; // {



endclass // }

`endif
