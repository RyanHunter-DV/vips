`ifndef Axi4MasterDriver__svh
`define Axi4MasterDriver__svh
`endif