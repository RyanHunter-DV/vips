`ifndef Axi4Vip__svh
`define Axi4Vip__svh
`endif
