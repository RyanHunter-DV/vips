`ifndef rhGpvDefines__svh
`define rhGpvDefines__svh
	`define RHGPV_MAX_VECTOR_WIDTH 1024
	`define RHGPV_MAX_CLOCK_WIDTH 16
	`define RHGPV_MAX_RESET_WIDTH 16
`endif
