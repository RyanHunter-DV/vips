package masterEnv;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "rhuMacros.svh"
	import rhudbg::*;

	import RhAhb5Vip::*;
	`include "masterEnv.svh"

endpackage
