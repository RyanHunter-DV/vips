`ifndef rhAhb5Vip__svh
`define rhAhb5Vip__svh

class RhAhb5Vip extends uvm_env;

	RhAhb5MstAgent   mst;
	RhAhb5SlvAgent   slv;
	RhAhb5ConfigBase config;
	RhuDebugger debug;

	`uvm_component_utils_begin(RhAhb5Vip)
	`uvm_component_utils_end
	function new(string name="RhAhb5Vip",uvm_component parent=null); // ##{{{
		super.new(name,parent);
		debug = new(this,"component");
	endfunction // ##}}}
	extern virtual function void build_phase(uvm_phase phase);
	extern function RhAhb5ConfigBase createConfig(RhAhb5MS_t m, string ifpath);
endclass
function void RhAhb5Vip::build_phase(uvm_phase phase);
	// This method is auto generated by cmd:Func
	if (config.isMaster()) begin
		mst = RhAhb5MstAgent::type_id::create("mst",this);
		mst.debug = debug;
		$cast(mst.config,config);
	end else begin
		slv = RhAhb5SlvAgent::type_id::create("slv",this);
		slv.debug = debug;
		$cast(slv.config,config);
	end
	debug.updateChildren(this);
endfunction
function RhAhb5ConfigBase RhAhb5Vip::createConfig(RhAhb5MS_t m, string ifpath);
	// This method is auto generated by cmd:Func
	// usage to set config:
	// config.setActivePassive(UVM_ACTIVE)
	// config.setMasterSlave(RHAHB5_MASTER)

	if (m==RHAHB5_MASTER) config = RhAhb5MstConfig::type_id::create("config");
	else config = RhAhb5SlvConfig::type_id::create("config");

	config.setMasterSlave(m);
	`debug($sformatf("calling getInterface with path: %s",ifpath))
	config.getInterface(ifpath);

	return config;
endfunction

`endif
