`ifndef Axi4SeqItem__svh
`define Axi4SeqItem__svh
`endif