`ifndef rhAhb5SlvMonitor__svh
`define rhAhb5SlvMonitor__svh

class RhAhb5SlvMonitor #(type REQ=uvm_sequence_item,RSP=REQ) extends RhMonitorBase;

	// request control phase port
	uvm_analysis_port#(REQ) reqCtrlP;
	// request data phase port, only available for write data
	uvm_analysis_port#(REQ) reqDataP;

	// response info, for read request, contains:
	// - data, resp, exokay
	// for write:
	// - resp, exokay
	uvm_analysis_port#(RSP) rspP;

	int outstandings= 0;
	RhAhb5SlvConfig config;
	// RhAhb5ReqTrans lastTr;
	uvm_event#(RhAhb5ReqTrans) writeReqEvent;
	uvm_event#(RhAhb5ReqTrans) reqEvent;

	`uvm_component_utils(RhAhb5SlvMonitor#(REQ,RSP))

	function new(string name="RhAhb5SlvMonitor",uvm_component parent=null);
		super.new(name,parent);
	endfunction

	// phases ##{{{
	extern function void build_phase (uvm_phase phase);
	extern function void connect_phase (uvm_phase phase);
	extern task run_phase (uvm_phase phase);
	// ##}}}

	// method group: main process ##{{{
	extern virtual task mainProcess();
	// ##}}}
	// method group: request monitor ##{{{
	extern task reqCtrlMonitor();
	extern task reqDataMonitor();
	// ##}}}

	// method group: response monitor ##{{{
	extern task rspMonitor();
	// ##}}}

	extern virtual task waitResetStateChanged(input RhResetState_enum c,output RhResetState_enum s);
endclass



//-----------------------CLASS BODY-----------------------//

task RhAhb5SlvMonitor::waitResetStateChanged(input RhResetState_enum c,output RhResetState_enum s);
	logic sig = logic'(c);
	config.getResetChanged(sig);
	s = RhResetState_enum'(sig);
endtask
task RhAhb5SlvMonitor::reqCtrlMonitor(); // ##{{{
	// This method is auto generated by cmd:Func
	// one execution of this task is monitoring one htrans request and send
	// through reqCtrlP
	logic [1:0] htrans;
	config.ifCtrl.clock();
	if (outstandings) begin
		while (config.ifCtrl.HREADY()!==1'b1) config.ifCtrl.clock(1);
	end
	htrans = config.ifCtrl.HTRANS();
	while (htrans!==1&&htrans!==2&&htrans!==3) begin
		config.ifCtrl.clock();
		htrans = config.ifCtrl.HTRANS();
	end
	if (htrans===1 || htrans===2 || htrans===3) begin
		RhAhb5ReqTrans req=new("reqCtrlTr");
		req.burst = config.ifCtrl.HBURST();
		req.addr  = config.ifCtrl.HADDR();
		req.prot  = config.ifCtrl.HPROT();
		req.lock  = config.ifCtrl.HMASTLOCK();
		req.trans = config.ifCtrl.HTRANS();
		req.size  = config.ifCtrl.HSIZE();
		req.nonsec= config.ifCtrl.HNONSEC();
		req.excl  = config.ifCtrl.HEXCL();
		req.write = config.ifCtrl.HWRITE();
		req.master= config.ifCtrl.HMASTER();
		req.stime = $time;
		if (req.write===1'b1) `rhudbgCall("write request detected, trigger writeReqEvent",writeReqEvent.trigger(req))
		`rhudbg($sformatf("collecting request by monitor:\n%s",req.sprint()))
		reqEvent.trigger(req); // for triggering rspMonitor
		req.etime =$time;
		reqCtrlP.write(req);
		`rhudbgCall($sformatf("do outstandings increment, current value(%0d)",outstandings),outstandings++)
	end
endtask // ##}}}
task RhAhb5SlvMonitor::reqDataMonitor(); // ##{{{
	// This method is auto generated by cmd:Func
	RhAhb5ReqTrans lastTr,req;
	writeReqEvent.wait_on();
	lastTr = writeReqEvent.get_trigger_data();
	writeReqEvent.reset();
	config.ifCtrl.clock();
	while (config.ifCtrl.HREADY()!=='b1) `rhudbgCall("waiting for HREADY=>1",config.ifCtrl.clock(1))
	req = new("reqDataTr");
	req.copy(lastTr);
	req.wdata = config.ifCtrl.HWDATA();
	`rhudbg($sformatf("collecting full write request transaction, with wdata:\n%s",req.sprint()))
	req.etime = $time; // flush etime
	reqDataP.write(req);
	// `rhudbgCall($sformatf("outstandings decrement, current value(%0d)",outstandings),outstandings--)
endtask // ##}}}
task RhAhb5SlvMonitor::rspMonitor(); // ##{{{
	// This method is auto generated by cmd:Func
	RhAhb5ReqTrans lastTr;
	RhAhb5RspTrans rsp;
	reqEvent.wait_on();
	lastTr = reqEvent.get_trigger_data();
	reqEvent.reset();
	`rhudbg($sformatf("reqEvent triggered, get req trans:\n%s",lastTr.sprint()))
	config.ifCtrl.clock();
	while (config.ifCtrl.HREADY()!== 1'b1)
		`rhudbgCall("in rspMonitor, waiting HREADY=>1",config.ifCtrl.clock(1))
	rsp = new("rspTr");
	rsp.stime = $time;
	rsp.iswrite = lastTr.write;
	rsp.exokay  = config.ifCtrl.HEXOKAY();
	rsp.resp    = config.ifCtrl.HRESP();
	if (lastTr.write===1'b0) rsp.rdata = config.ifCtrl.HRDATA();
	`rhudbg($sformatf("collecting response transaction:\n%s",rsp.sprint()))
	rsp.etime = $time;
	rspP.write(rsp);
	`rhudbgCall($sformatf("outstandings current value(%0d), decreasing to(%0d)",outstandings,outstandings-1),outstandings--)
endtask // ##}}}
task RhAhb5SlvMonitor::mainProcess(); // ##{{{
	// This method is auto generated by cmd:Func
	fork
		forever `rhudbgCall("starting reqCtrlMonitor ...",reqCtrlMonitor())
		forever `rhudbgCall("starting reqDataMonitor ...",reqDataMonitor())
		forever `rhudbgCall("starting rspMonitor ...",rspMonitor())
	join
endtask // ##}}}

function void RhAhb5SlvMonitor::build_phase(uvm_phase phase); // ##{{{
	super.build_phase(phase);
	reqCtrlP = new("reqCtrlP",this);
	reqDataP = new("reqDataP",this);
	rspP     = new("rspP",this);
	reqEvent = new("re");
	writeReqEvent = new("wre");
endfunction // ##}}}
function void RhAhb5SlvMonitor::connect_phase(uvm_phase phase); // ##{{{
	super.connect_phase(phase);
endfunction // ##}}}
task RhAhb5SlvMonitor::run_phase(uvm_phase phase); // ##{{{
	super.run_phase(phase);
endtask // ##}}}

`endif
