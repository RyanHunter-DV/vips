`ifndef Axi4MonitorBase__svh
`define Axi4MonitorBase__svh
`endif