class masterEnv extends uvm_env;



endclass
