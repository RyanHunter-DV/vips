`ifndef Axi4ResponseSeq__svh
`define Axi4ResponseSeq__svh
`endif