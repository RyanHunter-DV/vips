`ifndef Axi4MasterMonitor__svh
`define Axi4MasterMonitor__svh
`endif