package testsPkg;
	`include "uvm_macros.svh"
	`include "omosTestPkg.sv"

	import uvm_pkg::*;


	
endpackage
