`ifndef Axi4DriverBase__svh
`define Axi4DriverBase__svh
`endif