`ifndef Axi4BaseSeq__svh
`define Axi4BaseSeq__svh
`endif