`ifndef rhGpvTypes__svh
`define rhGpvTypes__svh



typedef bit [`RHGPV_MAX_VECTOR_WIDTH-1:0] bitVector_t;
typedef logic [`RHGPV_MAX_VECTOR_WIDTH-1:0] logicVector_t;




`endif
