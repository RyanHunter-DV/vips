`ifndef Axi4SlaveSeqr__svh
`define Axi4SlaveSeqr__svh
`endif