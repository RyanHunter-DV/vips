`ifndef rhAhb5Vip__svh
`define rhAhb5Vip__svh

class RhAhb5Vip extends uvm_env;

	parameter type REQ=RhAhb5ReqTrans;
	parameter type RSP=RhAhb5RspTrans;

	RhAhb5MstAgent#(REQ,RSP)   mst;
	RhAhb5SlvAgent#(REQ,RSP)   slv;
	RhAhb5ConfigBase config;
	RhuDebugger debug;
	RhAhb5MstSeqr seqr;

	uvm_analysis_export #(REQ) reqCtrlP;
	uvm_analysis_export #(REQ) reqDataP;
	uvm_analysis_export #(RSP) rspP;

	`uvm_component_utils_begin(RhAhb5Vip)
		`uvm_field_object(mst,UVM_ALL_ON)
		`uvm_field_object(slv,UVM_ALL_ON)
	`uvm_component_utils_end
	function new(string name="RhAhb5Vip",uvm_component parent=null); // ##{{{
		super.new(name,parent);
		debug = new(this,"component");
	endfunction // ##}}}
	// phases ##{{{
	// method group: build phase ##{{{
	extern virtual function void build_phase(uvm_phase phase);
	extern function void __localFieldsInitial__ ();
	// ##}}}
	extern function void connect_phase(uvm_phase phase);
	// ##}}}

	extern function RhAhb5ConfigBase createConfig(RhAhb5MS_t m, string ifpath);
endclass
function void RhAhb5Vip::__localFieldsInitial__(); // ##{{{
	reqCtrlP = new("reqCtrlP",this);
	reqDataP = new("reqDataP",this);
	rspP     = new("rspP",this);
endfunction // ##}}}
function void RhAhb5Vip::connect_phase(uvm_phase phase); // ##{{{
	super.connect_phase(phase);
	if (config.isMaster()) begin
		`debug("current is master mode, internal connecting with master")
		mst.reqCtrlP.connect(reqCtrlP);
		mst.reqDataP.connect(reqDataP);
		mst.rspP.connect(rspP);
	end else begin
		`debug("current is slave mode, internal connecting with slave")
		slv.reqCtrlP.connect(reqCtrlP);
		slv.reqDataP.connect(reqDataP);
		slv.rspP.connect(rspP);
	end
endfunction // ##}}}
function void RhAhb5Vip::build_phase(uvm_phase phase);
	// This method is auto generated by cmd:Func
	if (config.isMaster()) begin
		mst = RhAhb5MstAgent#(REQ,RSP)::type_id::create("mst",this);
		mst.debug = debug;
		`debugCall("setting master sequencer from the master agent",seqr = mst.seqr)
		$cast(mst.config,config);
	end else begin
		slv = RhAhb5SlvAgent#(REQ,RSP)::type_id::create("slv",this);
		slv.debug = debug;
		$cast(slv.config,config);
	end
	`debugCall("in build_phase, to init local fields",__localFieldsInitial__)
	debug.updateChildren(this);
endfunction
function RhAhb5ConfigBase RhAhb5Vip::createConfig(RhAhb5MS_t m, string ifpath);
	// This method is auto generated by cmd:Func
	// usage to set config:
	// config.setActivePassive(UVM_ACTIVE)
	// config.setMasterSlave(RHAHB5_MASTER)

	if (m==RHAHB5_MASTER) config = RhAhb5MstConfig::type_id::create("config");
	else config = RhAhb5SlvConfig::type_id::create("config");

	config.setMasterSlave(m);
	`debug($sformatf("calling getInterface with path: %s",ifpath))
	config.getInterface(ifpath);

	return config;
endfunction

`endif
