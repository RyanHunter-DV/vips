`ifndef rhGpvConfig__svh
`define rhGpvConfig__svh

class RhGpvConfig extends uvm_object;

	RhGpvIfCtrl ifCtrl;
	bit resetFeature;

	`uvm_object_utils_begin(RhGpvConfig)
	`uvm_object_utils_end

	function new(string name="RhGpvConfig");
		super.new(name);
	endfunction


	extern function void getInterface(string ifpath);
	extern function void driveVector(int s,int e,logicVector_t vector);
	// the return value starts from position 0 to the max size
	extern task sync(int pos, int cycle=1);
	extern function logicVector_t getOutSignal (int s,int e);
	extern function logicVector_t getInSignal (int s,int e);
	extern function logic getReset(int s);
	extern function void enableReset ();
endclass
function logic RhGpvConfig::getReset(int s); // ##{{{
	return ifCtrl.vif.getReset(s);
endfunction // ##}}}
function void RhGpvConfig::enableReset(); // ##{{{
	this.resetFeature = 1;
endfunction // ##}}}
// This code generated by snippet: 'func', if has any issue, pls report to RyanHunter
function logicVector_t RhGpvConfig::getOutSignal(int s,int e);
	return ifCtrl.vif.getVectorOut(s,e);
endfunction
function logicVector_t RhGpvConfig::getInSignal(int s,int e); // ##{{{
	return ifCtrl.vif.getVectorIn(s,e);
endfunction // ##}}}

task RhGpvConfig::sync(int pos, int cycle);
	`uvm_info("sync",$sformatf("calling ifCtrl.vif.sync(%0d,%0d)",pos,cycle),UVM_DEBUG)
	ifCtrl.vif.sync(pos,cycle);
	`uvm_info("sync",$sformatf("ifCtrl.vif.sync(%0d,%0d) synced",pos,cycle),UVM_DEBUG)
endtask

function void RhGpvConfig::driveVector(int s,int e,logicVector_t vector);
	logic bits[];
	int size = e-s+1;
	bits = new[size];
	for (int pos=s;pos<=e;pos++) begin
		bits[pos-s] = vector[pos];
	end
	ifCtrl.vif.driveVector(s,bits);
endfunction

function void RhGpvConfig::getInterface(string ifpath);
	if (!uvm_config_db#(RhGpvIfCtrl)::get(null,"*",ifpath,ifCtrl))
		`uvm_fatal("NCFG",$sformatf("interface path(%s) not found",ifpath))
endfunction

`endif
