`ifndef Axi4SlaveMonitor__svh
`define Axi4SlaveMonitor__svh
`endif