package env_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import RhGpVip::*;

	`include "rwaccessProtocol.svh"
	`include "env.svh"


endpackage
