`ifndef rhAhb5ResponderBase__svh
`define rhAhb5ResponderBase__svh

class RhAhb5ResponderBase extends uvm_object;

	`uvm_object_utils_begin(RhAhb5ResponderBase)
	`uvm_object_utils_end

	function new(string name="RhAhb5ResponderBase");
		super.new(name);
	endfunction


endclass

`endif
