`ifndef rhAhb5SlvConfig__svh
`define rhAhb5SlvConfig__svh

class RhAhb5SlvConfig extends RhAhb5ConfigBase;

	RhAhb5Response_t respMode;

	int lowDurationMins[string];
	int lowDurationMaxs[string];
	int highDurationMins[string];
	int highDurationMaxs[string];

	`uvm_object_utils_begin(RhAhb5SlvConfig)
		`uvm_field_enum(RhAhb5Response_t,respMode,UVM_ALL_ON)
	`uvm_object_utils_end

	function new(string name="RhAhb5SlvConfig");
		super.new(name);
		__setupDefaults__;
	endfunction

	// set response mode
	extern function void response(RhAhb5Response_t v);
	extern function bit israndom();
	extern function int lowDurationMin (string name);
	extern function int lowDurationMax (string name);
	extern function int highDurationMin (string name);
	extern function int highDurationMax (string name);
	extern function void __setupDefaults__ ();
endclass
function void RhAhb5SlvConfig::__setupDefaults__(); // ##{{{
	lowDurationMins["HREADY"] = 0;lowDurationMaxs["HREADY"] = 100;
	highDurationMins["HREADY"] = 0;highDurationMaxs["HREADY"] = 100;
endfunction // ##}}}
function int RhAhb5SlvConfig::lowDurationMin(string name); // ##{{{
	if (!lowDurationMins.exists(name)) begin
		`uvm_error("CFGE",$sformatf("attempt to get lowDurationMin(%s), which not configured",name))
		return 0;
	end
	return lowDurationMins[name];
endfunction // ##}}}
function int RhAhb5SlvConfig::lowDurationMax(string name); // ##{{{
	if (!lowDurationMaxs.exists(name)) begin
		`uvm_error("CFGE",$sformatf("attempt to get lowDurationMax(%s), which not configured",name))
		return 0;
	end
	return lowDurationMaxs[name];
endfunction // ##}}}
function int RhAhb5SlvConfig::highDurationMin(string name); // ##{{{
	if (!highDurationMins.exists(name)) begin
		`uvm_error("CFGE",$sformatf("attempt to get highDurationMin(%s), which not configured",name))
		return 0;
	end
	return highDurationMins[name];
endfunction // ##}}}
function int RhAhb5SlvConfig::highDurationMax(string name); // ##{{{
	if (!highDurationMaxs.exists(name)) begin
		`uvm_error("CFGE",$sformatf("attempt to get highDurationMax(%s), which not configured",name))
		return 0;
	end
	return highDurationMaxs[name];
endfunction // ##}}}

function bit RhAhb5SlvConfig::israndom(); // ##{{{
	// This method is auto generated by cmd:Func
	return (respMode==RHAHB5_RANDOM);
endfunction // ##}}}
function void RhAhb5SlvConfig::response(RhAhb5Response_t v); // ##{{{
	// This method is auto generated by cmd:Func
	respMode = v;
endfunction // ##}}}

`endif
