`ifndef Axi4Config__svh
`define Axi4Config__svh
`endif