`define RH_AXI4_IF_PARAM AW=32,DW=32,IW=16
