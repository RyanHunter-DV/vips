`ifndef omosEnvPkg__sv
`define omosEnvPkg__sv
package omosEnvPkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import rhudbg::*;
	import RhAhb5Vip::*;

	`include "omosEnv.svh"
endpackage
`endif
