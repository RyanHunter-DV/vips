package test_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import env_pkg::*;

	`include "selfTestSeq.svh"
	`include "baseTest.svh"
endpackage