`ifndef Axi4SlaveDriver__svh
`define Axi4SlaveDriver__svh
`endif