`ifndef RHAxi4MstAgent__svh
`define RHAxi4MstAgent__svh

class RHAxi4MstAgent extends uvm_agent;

	function new(string name="RHAxi4MstAgent",uvm_component parent=null);
		super.new(name,parent);
	endfunction

	

endclass

`endif
