`ifndef Axi4ResponseHandlerBase__svh
`define Axi4ResponseHandlerBase__svh
`endif