`ifndef Axi4SlaveAgent__svh
`define Axi4SlaveAgent__svh
`endif