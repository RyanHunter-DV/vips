`ifndef rhAhb5SlvConfig__svh
`define rhAhb5SlvConfig__svh

class RhAhb5SlvConfig extends RhAhb5ConfigBase;

	RhAhb5Response_t respMode;

	`uvm_object_utils_begin(RhAhb5SlvConfig)
		`uvm_field_enum(RhAhb5Response_t,respMode,UVM_ALL_ON)
	`uvm_object_utils_end

	function new(string name="RhAhb5SlvConfig");
		super.new(name);
	endfunction

	// set response mode
	extern function void response(RhAhb5Response_t v);
	extern function bit israndom();
endclass
function bit RhAhb5SlvConfig::israndom(); // ##{{{
	// This method is auto generated by cmd:Func
	return (respMode==RHAHB5_RANDOM);
endfunction // ##}}}
function void RhAhb5SlvConfig::response(RhAhb5Response_t v); // ##{{{
	// This method is auto generated by cmd:Func
	respMode = v;
endfunction // ##}}}

`endif
