`ifndef RhQLpiTests__sv
`define RhQLpiTests__sv

package RhQLpiTests;

	import uvm_pkg::*;
	import RhQLpiEnv::*; // env has imported vip package.

	`include "RhQLpiTestBase.svh"


endpackage

`endif