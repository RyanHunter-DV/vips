`ifndef Axi4ConfigBase__svh
`define Axi4ConfigBase__svh
`endif