`ifndef Axi4ResponseHandler__svh
`define Axi4ResponseHandler__svh
`endif