package ChiVipPkg;
/* Description, ChiVipPkg, 
*/
	import uvm_pkg::*;
	`include "rhlib.svh"

	import RhVipBase::*;
	

	`include "ChiVipTypedef.svh"

	`include "ChiSnDriver.svh"
endpackage