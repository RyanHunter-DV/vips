package env_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "rwaccessProtocol.svh"
	`include "env.svh"


endpackage