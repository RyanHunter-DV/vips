`ifndef RhPLpi__sv
`define RhPLpi__sv
package RhPLpi;
/* Description, RhPLpi, 
*/
	import uvm_pkg::*;
	`include "rhlib.svh"
	
endpackage
`endif