package MasterTestPkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import RhAhb5Vip::*;
	import masterEnv::*;

	`include "masterBaseTest.svh"

endpackage
