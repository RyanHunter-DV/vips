`ifndef Axi4MasterSeqr__svh
`define Axi4MasterSeqr__svh
`endif