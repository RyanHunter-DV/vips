package masterEnv;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	import RhAhb5Vip::*;
	`include "masterEnv.svh"

endpackage
