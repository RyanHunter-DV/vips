`ifndef RHAxi4ConfigBase__svh
`define RHAxi4ConfigBase__svh



`endif
