`ifndef Axi4VipLocalConfig__svh
`define Axi4VipLocalConfig__svh
`endif