`ifndef Axi4Interface__sv
`define Axi4Interface__sv
`endif